`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:21:37 11/16/2018 
// Design Name: 
// Module Name:    subtractor4bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module subtractor4bit(
    input [3:0] A,
    input [3:0] B,
    input [3:0] Cin,
    output [3:0] Cout
    );


endmodule
